
//main:	addi $2,$0,20 //initialise $2 =20
//		addi $3,$0,30 //initialise $3 =30
//		addi $5,$2,0 //initialise $5 =20
//		bne $5,$0,end //if val($5)!=val($0) branch to ‘end’
//		add $5,$2,$3 //$5=$2+$3
//end:	sw $5, 20($0) //write address 20 =20

module bne0_tb;
	reg clk;
	reg reset;
	integer i;
	wire [31:0] writedata, dataadr;
	wire memwrite;
	// instantiate device to be tested
	bne0 dut(clk, reset, writedata, dataadr, memwrite);
	
	// initialize test
	initial
	begin
		reset <= 1; # 22; reset <= 0;
	end
		// generate clock to sequence tests
	always
	begin
		clk <= 1; # 5; clk <= 0; # 5;
	end
		// check results
	always @ (negedge clk)
	begin
		if (memwrite) begin
			$display("%h %h\n", writedata,dataadr);
			if (dataadr === 20 & writedata === 20) begin
				$display ("Simulation succeeded");
				$stop;
			end else if (dataadr !== 80) begin
				$display ("Failed hehe %h and %h",writedata,dataadr);
				$stop;
			end
		end
	end
endmodule